//===============
// verification
//===============

//===============
// Import Package
//===============
import uvm_pkg::*;
`include "uvm_cros.svh"

//===============
//Interface
//===============
interface uart_if (input clk);
  logic rst_n;
  logic [7:0] tx_data;
  logic tx_start;
  logic tx;
  logic busy;
endinterface


//====================
//Class item_sequence
//====================





//===================
//Class uvm_sequence
//===================



//===================
//Class uvm_sequencer
//===================



//================
//Class uvm_driver
//================




//=================
//Class uvm_monitor
//=================





//===============
//Class uvm_agent
//===============




//====================
//Class uvm_scoreboard
//====================




//===============
//Class uvm_env
//===============





//===============
//Class base test
//===============





//====================
//    TOP MODULE
//==================== 




